`define PAWN   3'd0
`define KNIGHT 3'd1
`define BISHOP 3'd2
`define ROOK   3'd3
`define QUEEN  3'd4
`define KING   3'd5
`define EMPTY  3'd7

`define WHITE  1'b0
`define BLACK  1'b1

`define SM_FV        3'b000
`define SM_FP        3'b001
`define SM_FA        3'b010
`define SM_IDLE      3'b100
`define SM_DAAA      3'b101
`define SM_W         3'b110
`define SM_WD        3'b111

`define MM_EAV_EAA   2'b00
`define MM_DV_EAA    2'b01
`define MM_DA        2'b10
`define MM_NO_CHANGE 2'b11
